module compression ()

endmodule
