module text_compressor(input [7:0] binary_byte, 
								input clk, 
								output reg [6:0] compressed_byte
								);
always @(posedge clk)begin

if (binary_byte==8'b00100010) 
		compressed_byte= 7'b0;//string_out= " ";
	else if (binary_byte==8'b00100001)
		compressed_byte= 7'd1;//string_out= "!";
	else if (binary_byte==8'b00100011)
		compressed_byte= 7'd2;//string_out= "#";	
	else if (binary_byte==8'b00100100)
		compressed_byte= 7'd3;//string_out= "$";
	else if (binary_byte==8'b00100101)
		compressed_byte= 7'd4;//string_out= "%";
	else if (binary_byte==8'b00100110)
		compressed_byte= 7'd5;//string_out= "&";
	else if (binary_byte==8'b00100111)
		compressed_byte= 7'd6;//string_out= "'";
	else if (binary_byte==8'b00101000)
		compressed_byte= 7'd7;//string_out= "(";
	else if (binary_byte==8'b00101001)
		compressed_byte= 7'd8;//string_out= ")";
	else if (binary_byte==8'b00101010)
		compressed_byte= 7'd9;//string_out= "*";
	else if (binary_byte==8'b00101011)
		compressed_byte= 7'd10;//string_out= "+";
	else if (binary_byte==8'b00101100)
		compressed_byte= 7'd11;//string_out= ",";
	else if (binary_byte==8'b00101101)
		compressed_byte= 7'd12;//string_out= "-";	
	else if (binary_byte==8'b00101110)
		compressed_byte= 7'd13;//string_out= ".";
	else if (binary_byte==8'b00101111)
		compressed_byte= 7'd14;//string_out= "/";
	else if (binary_byte==8'b00110000)
		compressed_byte= 7'd15;//string_out= "0";
	else if (binary_byte==8'b00110001)
		compressed_byte= 7'd16;//string_out= "1";
	else if (binary_byte==8'b00110010)
		compressed_byte= 7'd17;//string_out= "2";
	else if (binary_byte==8'b00110011)
		compressed_byte= 7'd18;//string_out= "3";
	else if (binary_byte==8'b00110100)
		compressed_byte= 7'd19;//string_out= "4";
	else if (binary_byte==8'b00110101)
		compressed_byte= 7'd20;//string_out= "5";
	else if (binary_byte==8'b00110110)
		compressed_byte= 7'd21;//string_out= "6";
	else if (binary_byte==8'b00110111)
		compressed_byte= 7'd22;//string_out= "7";
	else if (binary_byte==8'b00111000)
		compressed_byte= 7'd23;//string_out= "8";
	else if (binary_byte==8'b00111001)
		compressed_byte= 7'd24;//string_out= "9";
	else if (binary_byte==8'b00111010)
		compressed_byte= 7'd25;//string_out= ":";
	else if (binary_byte==8'b00111011)
		compressed_byte= 7'd26;//string_out= ";";
	else if (binary_byte==8'b00111100)
		compressed_byte= 7'd27;//string_out= "<";
	else if (binary_byte==8'b00111101)
		compressed_byte= 7'd28;//string_out= "=";
	else if (binary_byte==8'b00111110)
		compressed_byte= 7'd29;//string_out= ">";
	else if (binary_byte==8'b00111111)
		compressed_byte= 7'd30;//string_out= "?";
	else if (binary_byte==8'b01000000)
		compressed_byte= 7'd31;//string_out= "@";
	else if (binary_byte==8'b01000001)
		compressed_byte= 7'd32;//string_out= "A";
	else if (binary_byte==8'b01000010)
		compressed_byte= 7'd33;//string_out= "B";
	else if (binary_byte==8'b01000011)
		compressed_byte= 7'd34;//string_out= "C";
	else if (binary_byte==8'b01000100)
		compressed_byte= 7'd35;//string_out= "D";
	else if (binary_byte==8'b01000101)
		compressed_byte= 7'd36;//string_out= "E";
	else if (binary_byte==8'b01000110)
		compressed_byte= 7'd37;//string_out= "F";
	else if (binary_byte==8'b01000111)
		compressed_byte= 7'd38;//string_out= "G";
	else if (binary_byte==8'b01001000)
		compressed_byte= 7'd39;//string_out= "H";
	else if (binary_byte==8'b01001001)
		compressed_byte= 7'd40;//string_out= "I";
	else if (binary_byte==8'b01001010)
		compressed_byte= 7'd41;//string_out= "J";
	else if (binary_byte==8'b01001011)
		compressed_byte= 7'd42;//string_out= "K";
	else if (binary_byte==8'b01001100)
		compressed_byte= 7'd43;//string_out= "L";
	else if (binary_byte==8'b01001101)
		compressed_byte= 7'd44;//string_out= "M";
	else if (binary_byte==8'b01001110)
		compressed_byte= 7'd45;//string_out= "N";
	else if (binary_byte==8'b01001111)
		compressed_byte= 7'd46;//string_out= "O";
	else if (binary_byte==8'b01010000)
		compressed_byte= 7'd47;//string_out= "P";
	else if (binary_byte==8'b01010001)
		compressed_byte= 7'd48;//string_out= "Q";
	else if (binary_byte==8'b01010010)
		compressed_byte= 7'd49;//string_out= "R";
	else if (binary_byte==8'b01010011)
		compressed_byte= 7'd50;//string_out= "S";
	else if (binary_byte==8'b01010100)
		compressed_byte= 7'd51;//string_out= "T";
	else if (binary_byte==8'b01010101)
		compressed_byte= 7'd52;//string_out= "U";
	else if (binary_byte==8'b01010110)
		compressed_byte= 7'd53;//string_out= "V";
	else if (binary_byte==8'b01010111)
		compressed_byte= 7'd54;//string_out= "W";	
	else if (binary_byte==8'b01010000)
		compressed_byte= 7'd55;//string_out= "X";
	else if (binary_byte==8'b01011001)
		compressed_byte= 7'd56;//string_out= "Y";
	else if (binary_byte==8'b01011010)
		compressed_byte= 7'd57;//string_out= "Z";
	else if (binary_byte==8'b01011011)
		compressed_byte= 7'd58;//string_out= "[";
	else if (binary_byte==8'b01011100)
		compressed_byte= 7'd59;//string_out= "";//\
	else if (binary_byte==8'b01011101)
		compressed_byte= 7'd60;//string_out= "]";
	else if (binary_byte==8'b01011110)
		compressed_byte= 7'd61;//string_out= "^";
	else if (binary_byte==8'b01011111)
		compressed_byte= 7'd62;//string_out= "_";
	else if (binary_byte==8'b01100000)
		compressed_byte= 7'd63;//string_out= "`";
	else if (binary_byte==8'b01100001)
		compressed_byte= 7'd64;//string_out= "a";
	else if (binary_byte==8'b01100010)
		compressed_byte= 7'd65;//string_out= "b";
	else if (binary_byte==8'b01100011)
		compressed_byte= 7'd66;//string_out= "c";
	else if (binary_byte==8'b01100100)
		compressed_byte= 7'd67;//string_out= "d";
	else if (binary_byte==8'b01100101)
		compressed_byte= 7'd68;//string_out= "e";
	else if (binary_byte==8'b01100110)
		compressed_byte= 7'd69;//string_out= "f";
	else if (binary_byte==8'b01100111)
		compressed_byte= 7'd70;//string_out= "g";
	else if (binary_byte==8'b01101000)
		compressed_byte= 7'd71;//string_out= "h";
	else if (binary_byte==8'b01101001)
		compressed_byte= 7'd72;//string_out= "i";
	else if (binary_byte==8'b01101010)
		compressed_byte= 7'd73;//string_out= "j";
	else if (binary_byte==8'b01101011)
		compressed_byte= 7'd74;//string_out= "k";
	else if (binary_byte==8'b01101100)
		compressed_byte= 7'd75;//string_out= "l";
	else if (binary_byte==8'b01101101)
		compressed_byte= 7'd76;//string_out= "m";
	else if (binary_byte==8'b01101110)
		compressed_byte= 7'd77;//string_out= "n";
	else if (binary_byte==8'b01101111)
		compressed_byte= 7'd78;//string_out= "o";
	else if (binary_byte==8'b01110000)
		compressed_byte= 7'd79;//string_out= "p";
	else if (binary_byte==8'b01110001)
		compressed_byte= 7'd80;//string_out= "q";
	else if (binary_byte==8'b01110010)
		compressed_byte= 7'd81;//string_out= "r";
	else if (binary_byte==8'b01110011)
		compressed_byte= 7'd82;//string_out= "s";
	else if (binary_byte==8'b01110100)
		compressed_byte= 7'd83;//string_out= "t";
	else if (binary_byte==8'b01110101)
		compressed_byte= 7'd84;//string_out= "u";
	else if (binary_byte==8'b01110110)
		compressed_byte= 7'd85;//string_out= "v";	
	else if (binary_byte==8'b01110111)
		compressed_byte= 7'd86;//string_out= "w";
	else if (binary_byte==8'b01111000)
		compressed_byte= 7'd87;//string_out= "x";
	else if (binary_byte==8'b01111001)
		compressed_byte= 7'd88;//string_out= "y";
	else if (binary_byte==8'b01111010)
		compressed_byte= 7'd89;//string_out= "z";
	else if (binary_byte==8'b01111011)
		compressed_byte= 7'd90;//string_out= "{";
	else if (binary_byte==8'b01111100)
		compressed_byte= 7'd91;//string_out= "|";
	else if (binary_byte==8'b01111101)
		compressed_byte= 7'd92;//string_out= "}";
	else if (binary_byte==8'b01111111)
		compressed_byte=7'd93;//string out="DEL"
	else if (binary_byte==8'b10000000)
		compressed_byte=7'd94;//string_out="NUL"
	else compressed_byte= 7'd95;//string_out="~";
	
end

endmodule